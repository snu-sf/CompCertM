Require Import AST Coqlib.
Require Import Asm.
Require Import sflib.
Require Import AsmC Mod.
Require Import Header.

Definition lb0: label := 1%positive.
Definition code: list instruction :=
  [
    Ptestq_rr RDI RDI ;
      Pjcc Cond_s lb0 ;
      Pxorpd_f XMM0 ;
      (* note: actual code is pxor, but it it prints xorpd *)
      (* it also prints the same thing: Pxorps_f XMM0 ; *)
      Pcvtsl2ss_fr XMM0 RDI ;
      Pret ;

      Plabel lb0 ;
      Pmov_rr RAX RDI ;
      Pshrq_ri RAX Integers.Int.one ;
      Pandq_ri RDI Integers.Int64.one ;
      Porq_rr RAX RDI ;
      Pxorpd_f XMM0 ;
      Pcvtsl2ss_fr XMM0 RAX ;
      Padds_ff XMM0 XMM0 ;
      Pret
  ].

Definition func: function :=
  mkfunction (mksignature [Tlong] (Some Tsingle) cc_default) code
.

Definition prog: program := mkprogram [(func_id, (Gfun (Internal func)))] [func_id ; main_id] main_id.

Definition md: Mod.t := AsmC.module prog.

Hint Unfold md prog func code.













Extract Inductive list => "list" [ "[]" "(::)" ].
Extract Inlined Constant Datatypes.fst => "fst".
Extract Inlined Constant Datatypes.snd => "snd".
Extract Inductive prod => "(*)"  [ "(,)" ].
(* Recursive Extraction utof_program. *)
Extraction lb0.
Extraction code.
Extraction func.
Extraction func_id.
Extraction prog.


(****************************** ORIGINAL *****************************************)
(* FUNCTION(__compcert_i64_utof) *)
(*         testq   %rdi, %rdi *)
(*         js      1f *)
(*         pxor    %xmm0, %xmm0            // if < 2^63, *)
(*         cvtsi2ssq %rdi, %xmm0           // convert as if signed *)
(*         ret *)
(* 1:                                      // if >= 2^63, use round-to-odd trick *)
(*         movq    %rdi, %rax *)
(*         shrq    %rax *)
(*         andq    $1, %rdi *)
(*         orq     %rdi, %rax              // (arg >> 1) | (arg & 1) *)
(*         pxor    %xmm0, %xmm0 *)
(*         cvtsi2ssq %rax, %xmm0           // convert as if signed *)
(*         addss   %xmm0, %xmm0            // multiply result by 2.0 *)
(*         ret *)
(* ENDFUNCTION(__compcert_i64_utof) *)




(****************************** FROM COQ *****************************************)
(* # File generated by CompCert 3.4 *)
(* # Command line: --help *)
(*         .text *)
(*         .align  16 *)
(*         .globl $2 *)
(* $2: *)
(*         .cfi_startproc *)
(*         testq   %rdi, %rdi *)
(*         jmp     .L100 *)
(*         xorpd   %xmm0, %xmm0 *)
(*         cvtsi2ssq %rdi, %xmm0 *)
(*         ret *)
(* .L100: *)
(*         movq    %rdi, %rax *)
(*         shrq    $1, %rax *)
(*         andq    $1, %rdi *)
(*         orq     %rdi, %rax *)
(*         xorpd   %xmm0, %xmm0 *)
(*         cvtsi2ssq %rax, %xmm0 *)
(*         addss   %xmm0, %xmm0 *)
(*         ret *)
(*         .cfi_endproc *)
(*         .type   $2, @function *)
(*         .size   $2, . - $2 *)